library verilog;
use verilog.vl_types.all;
entity circuiteria_vlg_vec_tst is
end circuiteria_vlg_vec_tst;
