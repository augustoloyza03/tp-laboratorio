library verilog;
use verilog.vl_types.all;
entity parteD_vlg_vec_tst is
end parteD_vlg_vec_tst;
