library verilog;
use verilog.vl_types.all;
entity circuiteria_vlg_check_tst is
    port(
        finDATO         : in     vl_logic;
        finDIR          : in     vl_logic;
        soy             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end circuiteria_vlg_check_tst;
