library verilog;
use verilog.vl_types.all;
entity parteB_vlg_vec_tst is
end parteB_vlg_vec_tst;
