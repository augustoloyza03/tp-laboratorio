library verilog;
use verilog.vl_types.all;
entity parteD_vlg_check_tst is
    port(
        Z0              : in     vl_logic;
        Z1              : in     vl_logic;
        Z2              : in     vl_logic;
        Z3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end parteD_vlg_check_tst;
