library verilog;
use verilog.vl_types.all;
entity Block1_vlg_check_tst is
    port(
        Bout            : in     vl_logic;
        Z0              : in     vl_logic;
        Z1              : in     vl_logic;
        Z2              : in     vl_logic;
        Z3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Block1_vlg_check_tst;
